// Copyright 2022 ETH Zurich and University of Bologna.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51
//
// Fabian Schuiki <fschuiki@iis.ee.ethz.ch>
// Florian Zaruba <zarubaf@iis.ee.ethz.ch>
// Stefan Mach <smach@iis.ee.ethz.ch>
// Thomas Benz <tbenz@iis.ee.ethz.ch>
// Paul Scheffler <paulsc@iis.ee.ethz.ch>
// Wolfgang Roenninger <wroennin@iis.ee.ethz.ch>
//
// AUTOMATICALLY GENERATED by bin2sv.py; edit the script instead.

module bootrom #(
    parameter int unsigned AddrWidth = 32,
    parameter int unsigned DataWidth = 32
)(
    input  logic                 clk_i,
    input  logic                 rst_ni,
    input  logic                 req_i,
    input  logic [AddrWidth-1:0] addr_i,
    output logic [DataWidth-1:0] data_o
);
    localparam unsigned NumWords = 1024;
    logic [$clog2(NumWords)-1:0] word;

    assign word = addr_i / (DataWidth / 8);

    always_comb begin
        data_o = '0;
        unique case (word)
        000: data_o = 32'h301022f3 /* 0x0000 */;
            001: data_o = 32'h0202ce63 /* 0x0004 */;
            002: data_o = 32'hf1402573 /* 0x0008 */;
            003: data_o = 32'h6f000297 /* 0x000c */;
            004: data_o = 32'hffc2b283 /* 0x0010 */;
            005: data_o = 32'h30529073 /* 0x0014 */;
            006: data_o = 32'h30046073 /* 0x0018 */;
            007: data_o = 32'h000802b7 /* 0x001c */;
            008: data_o = 32'h00828293 /* 0x0020 */;
            009: data_o = 32'h30429073 /* 0x0024 */;
            010: data_o = 32'h10500073 /* 0x0028 */;
            011: data_o = 32'h6f000297 /* 0x002c */;
            012: data_o = 32'hffc2b283 /* 0x0030 */;
            013: data_o = 32'h0002a283 /* 0x0034 */;
            014: data_o = 32'h000280e7 /* 0x0038 */;
            015: data_o = 32'hfcdff06f /* 0x003c */;
            016: data_o = 32'hf1502473 /* 0x0040 */;
            017: data_o = 32'h02841413 /* 0x0044 */;
            018: data_o = 32'h6f000197 /* 0x0048 */;
            019: data_o = 32'hfd01b183 /* 0x004c */;
            020: data_o = 32'h0081f1b3 /* 0x0050 */;
            021: data_o = 32'h6f000117 /* 0x0054 */;
            022: data_o = 32'hfcc13103 /* 0x0058 */;
            023: data_o = 32'h00817133 /* 0x005c */;
            024: data_o = 32'h6f000317 /* 0x0060 */;
            025: data_o = 32'hfb033303 /* 0x0064 */;
            026: data_o = 32'h30531073 /* 0x0068 */;
            027: data_o = 32'h464000ef /* 0x006c */;
            028: data_o = 32'h0010029b /* 0x0070 */;
            029: data_o = 32'h01f29293 /* 0x0074 */;
            030: data_o = 32'h000280e7 /* 0x0078 */;
            031: data_o = 32'hf85ff06f /* 0x007c */;
            032: data_o = 32'h10500073 /* 0x0080 */;
            033: data_o = 32'hffdff06f /* 0x0084 */;
            034: data_o = 32'hff010113 /* 0x0088 */;
            035: data_o = 32'h00813423 /* 0x008c */;
            036: data_o = 32'h01002717 /* 0x0090 */;
            037: data_o = 32'hf8470713 /* 0x0094 */;
            038: data_o = 32'h01010413 /* 0x0098 */;
            039: data_o = 32'h00a76733 /* 0x009c */;
            040: data_o = 32'h00074783 /* 0x00a0 */;
            041: data_o = 32'h0207f793 /* 0x00a4 */;
            042: data_o = 32'hfe078ce3 /* 0x00a8 */;
            043: data_o = 32'h01002797 /* 0x00ac */;
            044: data_o = 32'hf5478793 /* 0x00b0 */;
            045: data_o = 32'h00f56533 /* 0x00b4 */;
            046: data_o = 32'h00b50023 /* 0x00b8 */;
            047: data_o = 32'h00813403 /* 0x00bc */;
            048: data_o = 32'h01010113 /* 0x00c0 */;
            049: data_o = 32'h00008067 /* 0x00c4 */;
            050: data_o = 32'hff010113 /* 0x00c8 */;
            051: data_o = 32'h00813423 /* 0x00cc */;
            052: data_o = 32'h01002717 /* 0x00d0 */;
            053: data_o = 32'hf4470713 /* 0x00d4 */;
            054: data_o = 32'h01010413 /* 0x00d8 */;
            055: data_o = 32'h00a76733 /* 0x00dc */;
            056: data_o = 32'h00074783 /* 0x00e0 */;
            057: data_o = 32'h0017f793 /* 0x00e4 */;
            058: data_o = 32'hfe078ce3 /* 0x00e8 */;
            059: data_o = 32'h00813403 /* 0x00ec */;
            060: data_o = 32'h01002797 /* 0x00f0 */;
            061: data_o = 32'hf1078793 /* 0x00f4 */;
            062: data_o = 32'h00f56533 /* 0x00f8 */;
            063: data_o = 32'h00054503 /* 0x00fc */;
            064: data_o = 32'h01010113 /* 0x0100 */;
            065: data_o = 32'h00008067 /* 0x0104 */;
            066: data_o = 32'hfe010113 /* 0x0108 */;
            067: data_o = 32'h00813823 /* 0x010c */;
            068: data_o = 32'h00913423 /* 0x0110 */;
            069: data_o = 32'h01213023 /* 0x0114 */;
            070: data_o = 32'h00113c23 /* 0x0118 */;
            071: data_o = 32'h02010413 /* 0x011c */;
            072: data_o = 32'h00050913 /* 0x0120 */;
            073: data_o = 32'h00058493 /* 0x0124 */;
            074: data_o = 32'h0004c583 /* 0x0128 */;
            075: data_o = 32'h02059a63 /* 0x012c */;
            076: data_o = 32'h01002517 /* 0x0130 */;
            077: data_o = 32'hee450513 /* 0x0134 */;
            078: data_o = 32'h01256533 /* 0x0138 */;
            079: data_o = 32'h00054783 /* 0x013c */;
            080: data_o = 32'h0407f793 /* 0x0140 */;
            081: data_o = 32'hfe078ce3 /* 0x0144 */;
            082: data_o = 32'h01813083 /* 0x0148 */;
            083: data_o = 32'h01013403 /* 0x014c */;
            084: data_o = 32'h00813483 /* 0x0150 */;
            085: data_o = 32'h00013903 /* 0x0154 */;
            086: data_o = 32'h02010113 /* 0x0158 */;
            087: data_o = 32'h00008067 /* 0x015c */;
            088: data_o = 32'h00090513 /* 0x0160 */;
            089: data_o = 32'hf25ff0ef /* 0x0164 */;
            090: data_o = 32'h00148493 /* 0x0168 */;
            091: data_o = 32'hfbdff06f /* 0x016c */;
            092: data_o = 32'hfa010113 /* 0x0170 */;
            093: data_o = 32'h04813823 /* 0x0174 */;
            094: data_o = 32'h05213023 /* 0x0178 */;
            095: data_o = 32'h06010413 /* 0x017c */;
            096: data_o = 32'h03313c23 /* 0x0180 */;
            097: data_o = 32'h03413823 /* 0x0184 */;
            098: data_o = 32'h03513423 /* 0x0188 */;
            099: data_o = 32'h03613023 /* 0x018c */;
            100: data_o = 32'h04113c23 /* 0x0190 */;
            101: data_o = 32'h04913423 /* 0x0194 */;
            102: data_o = 32'h01713c23 /* 0x0198 */;
            103: data_o = 32'h00000797 /* 0x019c */;
            104: data_o = 32'h7e478793 /* 0x01a0 */;
            105: data_o = 32'h0007b783 /* 0x01a4 */;
            106: data_o = 32'h00050a13 /* 0x01a8 */;
            107: data_o = 32'h00058993 /* 0x01ac */;
            108: data_o = 32'hfaf43023 /* 0x01b0 */;
            109: data_o = 32'h00000797 /* 0x01b4 */;
            110: data_o = 32'h7d478793 /* 0x01b8 */;
            111: data_o = 32'h0007b783 /* 0x01bc */;
            112: data_o = 32'h00060a93 /* 0x01c0 */;
            113: data_o = 32'h00000913 /* 0x01c4 */;
            114: data_o = 32'hfaf43423 /* 0x01c8 */;
            115: data_o = 32'hffc00b13 /* 0x01cc */;
            116: data_o = 32'h00090b9b /* 0x01d0 */;
            117: data_o = 32'h053be263 /* 0x01d4 */;
            118: data_o = 32'h01002717 /* 0x01d8 */;
            119: data_o = 32'he3c70713 /* 0x01dc */;
            120: data_o = 32'h00074783 /* 0x01e0 */;
            121: data_o = 32'h0407f793 /* 0x01e4 */;
            122: data_o = 32'hfe078ce3 /* 0x01e8 */;
            123: data_o = 32'h05813083 /* 0x01ec */;
            124: data_o = 32'h05013403 /* 0x01f0 */;
            125: data_o = 32'h04813483 /* 0x01f4 */;
            126: data_o = 32'h04013903 /* 0x01f8 */;
            127: data_o = 32'h03813983 /* 0x01fc */;
            128: data_o = 32'h03013a03 /* 0x0200 */;
            129: data_o = 32'h02813a83 /* 0x0204 */;
            130: data_o = 32'h02013b03 /* 0x0208 */;
            131: data_o = 32'h01813b83 /* 0x020c */;
            132: data_o = 32'h06010113 /* 0x0210 */;
            133: data_o = 32'h00008067 /* 0x0214 */;
            134: data_o = 32'h00fbf793 /* 0x0218 */;
            135: data_o = 32'h06079063 /* 0x021c */;
            136: data_o = 32'h040a8e63 /* 0x0220 */;
            137: data_o = 32'h00d00593 /* 0x0224 */;
            138: data_o = 32'h00000513 /* 0x0228 */;
            139: data_o = 32'he5dff0ef /* 0x022c */;
            140: data_o = 32'h00a00593 /* 0x0230 */;
            141: data_o = 32'h00000513 /* 0x0234 */;
            142: data_o = 32'he51ff0ef /* 0x0238 */;
            143: data_o = 32'h01c00493 /* 0x023c */;
            144: data_o = 32'h009bd7bb /* 0x0240 */;
            145: data_o = 32'hfb040713 /* 0x0244 */;
            146: data_o = 32'h00f7f793 /* 0x0248 */;
            147: data_o = 32'h00f707b3 /* 0x024c */;
            148: data_o = 32'hff07c583 /* 0x0250 */;
            149: data_o = 32'h00000513 /* 0x0254 */;
            150: data_o = 32'hffc4849b /* 0x0258 */;
            151: data_o = 32'he2dff0ef /* 0x025c */;
            152: data_o = 32'hff6490e3 /* 0x0260 */;
            153: data_o = 32'h03a00593 /* 0x0264 */;
            154: data_o = 32'h00000513 /* 0x0268 */;
            155: data_o = 32'he1dff0ef /* 0x026c */;
            156: data_o = 32'h02000593 /* 0x0270 */;
            157: data_o = 32'h00000513 /* 0x0274 */;
            158: data_o = 32'he11ff0ef /* 0x0278 */;
            159: data_o = 32'h012a07b3 /* 0x027c */;
            160: data_o = 32'h0007c483 /* 0x0280 */;
            161: data_o = 32'hfb040713 /* 0x0284 */;
            162: data_o = 32'h00000513 /* 0x0288 */;
            163: data_o = 32'h0044d793 /* 0x028c */;
            164: data_o = 32'h00f707b3 /* 0x0290 */;
            165: data_o = 32'hff07c583 /* 0x0294 */;
            166: data_o = 32'h00f4f493 /* 0x0298 */;
            167: data_o = 32'h00190913 /* 0x029c */;
            168: data_o = 32'hde9ff0ef /* 0x02a0 */;
            169: data_o = 32'hfb040793 /* 0x02a4 */;
            170: data_o = 32'h009784b3 /* 0x02a8 */;
            171: data_o = 32'hff04c583 /* 0x02ac */;
            172: data_o = 32'h00000513 /* 0x02b0 */;
            173: data_o = 32'hdd5ff0ef /* 0x02b4 */;
            174: data_o = 32'h02000593 /* 0x02b8 */;
            175: data_o = 32'h00000513 /* 0x02bc */;
            176: data_o = 32'hdc9ff0ef /* 0x02c0 */;
            177: data_o = 32'hf0dff06f /* 0x02c4 */;
            178: data_o = 32'hff010113 /* 0x02c8 */;
            179: data_o = 32'h00813423 /* 0x02cc */;
            180: data_o = 32'h01010413 /* 0x02d0 */;
            181: data_o = 32'h00000713 /* 0x02d4 */;
            182: data_o = 32'h00000793 /* 0x02d8 */;
            183: data_o = 32'h0007069b /* 0x02dc */;
            184: data_o = 32'h00b6ea63 /* 0x02e0 */;
            185: data_o = 32'h00813403 /* 0x02e4 */;
            186: data_o = 32'h00078513 /* 0x02e8 */;
            187: data_o = 32'h01010113 /* 0x02ec */;
            188: data_o = 32'h00008067 /* 0x02f0 */;
            189: data_o = 32'h00e506b3 /* 0x02f4 */;
            190: data_o = 32'h0006c683 /* 0x02f8 */;
            191: data_o = 32'h00170713 /* 0x02fc */;
            192: data_o = 32'h00d787b3 /* 0x0300 */;
            193: data_o = 32'h0ff7f793 /* 0x0304 */;
            194: data_o = 32'hfd5ff06f /* 0x0308 */;
            195: data_o = 32'hff010113 /* 0x030c */;
            196: data_o = 32'h00813423 /* 0x0310 */;
            197: data_o = 32'h01010413 /* 0x0314 */;
            198: data_o = 32'h00000793 /* 0x0318 */;
            199: data_o = 32'h0007871b /* 0x031c */;
            200: data_o = 32'h00c76863 /* 0x0320 */;
            201: data_o = 32'h00813403 /* 0x0324 */;
            202: data_o = 32'h01010113 /* 0x0328 */;
            203: data_o = 32'h00008067 /* 0x032c */;
            204: data_o = 32'h00f58733 /* 0x0330 */;
            205: data_o = 32'h00074683 /* 0x0334 */;
            206: data_o = 32'h00f50733 /* 0x0338 */;
            207: data_o = 32'h00178793 /* 0x033c */;
            208: data_o = 32'h00d70023 /* 0x0340 */;
            209: data_o = 32'hfd9ff06f /* 0x0344 */;
            210: data_o = 32'hbb010113 /* 0x0348 */;
            211: data_o = 32'h44813023 /* 0x034c */;
            212: data_o = 32'h42913c23 /* 0x0350 */;
            213: data_o = 32'h43413023 /* 0x0354 */;
            214: data_o = 32'h41513c23 /* 0x0358 */;
            215: data_o = 32'h41613823 /* 0x035c */;
            216: data_o = 32'h41713423 /* 0x0360 */;
            217: data_o = 32'h44113423 /* 0x0364 */;
            218: data_o = 32'h43213823 /* 0x0368 */;
            219: data_o = 32'h43313423 /* 0x036c */;
            220: data_o = 32'h45010413 /* 0x0370 */;
            221: data_o = 32'h00058b93 /* 0x0374 */;
            222: data_o = 32'h01500593 /* 0x0378 */;
            223: data_o = 32'h00050493 /* 0x037c */;
            224: data_o = 32'h00000a13 /* 0x0380 */;
            225: data_o = 32'hd05ff0ef /* 0x0384 */;
            226: data_o = 32'h00400b13 /* 0x0388 */;
            227: data_o = 32'h00100a93 /* 0x038c */;
            228: data_o = 32'h00048513 /* 0x0390 */;
            229: data_o = 32'hd35ff0ef /* 0x0394 */;
            230: data_o = 32'h00050993 /* 0x0398 */;
            231: data_o = 32'h05651663 /* 0x039c */;
            232: data_o = 32'h00048513 /* 0x03a0 */;
            233: data_o = 32'h00600593 /* 0x03a4 */;
            234: data_o = 32'hce1ff0ef /* 0x03a8 */;
            235: data_o = 32'h00048513 /* 0x03ac */;
            236: data_o = 32'h00000597 /* 0x03b0 */;
            237: data_o = 32'h42058593 /* 0x03b4 */;
            238: data_o = 32'hd51ff0ef /* 0x03b8 */;
            239: data_o = 32'h44813083 /* 0x03bc */;
            240: data_o = 32'h44013403 /* 0x03c0 */;
            241: data_o = 32'h43813483 /* 0x03c4 */;
            242: data_o = 32'h43013903 /* 0x03c8 */;
            243: data_o = 32'h42813983 /* 0x03cc */;
            244: data_o = 32'h42013a03 /* 0x03d0 */;
            245: data_o = 32'h41813a83 /* 0x03d4 */;
            246: data_o = 32'h41013b03 /* 0x03d8 */;
            247: data_o = 32'h40813b83 /* 0x03dc */;
            248: data_o = 32'h45010113 /* 0x03e0 */;
            249: data_o = 32'h00008067 /* 0x03e4 */;
            250: data_o = 32'hfff9879b /* 0x03e8 */;
            251: data_o = 32'h0ff7f793 /* 0x03ec */;
            252: data_o = 32'h01800593 /* 0x03f0 */;
            253: data_o = 32'h0afae263 /* 0x03f4 */;
            254: data_o = 32'h00048513 /* 0x03f8 */;
            255: data_o = 32'hccdff0ef /* 0x03fc */;
            256: data_o = 32'h00050913 /* 0x0400 */;
            257: data_o = 32'h00048513 /* 0x0404 */;
            258: data_o = 32'hcc1ff0ef /* 0x0408 */;
            259: data_o = 32'hfff54513 /* 0x040c */;
            260: data_o = 32'h0ff57513 /* 0x0410 */;
            261: data_o = 32'h09251063 /* 0x0414 */;
            262: data_o = 32'h40000913 /* 0x0418 */;
            263: data_o = 32'h01599463 /* 0x041c */;
            264: data_o = 32'h08000913 /* 0x0420 */;
            265: data_o = 32'h00000993 /* 0x0424 */;
            266: data_o = 32'h0009879b /* 0x0428 */;
            267: data_o = 32'h00048513 /* 0x042c */;
            268: data_o = 32'h0527c663 /* 0x0430 */;
            269: data_o = 32'hc95ff0ef /* 0x0434 */;
            270: data_o = 32'h0009091b /* 0x0438 */;
            271: data_o = 32'h00050993 /* 0x043c */;
            272: data_o = 32'h00090593 /* 0x0440 */;
            273: data_o = 32'hbb040513 /* 0x0444 */;
            274: data_o = 32'he81ff0ef /* 0x0448 */;
            275: data_o = 32'h04a99463 /* 0x044c */;
            276: data_o = 32'h00600593 /* 0x0450 */;
            277: data_o = 32'h00048513 /* 0x0454 */;
            278: data_o = 32'hc31ff0ef /* 0x0458 */;
            279: data_o = 32'h020a1513 /* 0x045c */;
            280: data_o = 32'h02055513 /* 0x0460 */;
            281: data_o = 32'h00090613 /* 0x0464 */;
            282: data_o = 32'hbb040593 /* 0x0468 */;
            283: data_o = 32'h01750533 /* 0x046c */;
            284: data_o = 32'he9dff0ef /* 0x0470 */;
            285: data_o = 32'h01490a3b /* 0x0474 */;
            286: data_o = 32'hf19ff06f /* 0x0478 */;
            287: data_o = 32'hc4dff0ef /* 0x047c */;
            288: data_o = 32'hbb040793 /* 0x0480 */;
            289: data_o = 32'h013787b3 /* 0x0484 */;
            290: data_o = 32'h00a78023 /* 0x0488 */;
            291: data_o = 32'h00198993 /* 0x048c */;
            292: data_o = 32'hf99ff06f /* 0x0490 */;
            293: data_o = 32'h01500593 /* 0x0494 */;
            294: data_o = 32'h00048513 /* 0x0498 */;
            295: data_o = 32'hbedff0ef /* 0x049c */;
            296: data_o = 32'hef1ff06f /* 0x04a0 */;
            297: data_o = 32'hff010113 /* 0x04a4 */;
            298: data_o = 32'h00813423 /* 0x04a8 */;
            299: data_o = 32'h01010413 /* 0x04ac */;
            300: data_o = 32'hb00027f3 /* 0x04b0 */;
            301: data_o = 32'h00a787b3 /* 0x04b4 */;
            302: data_o = 32'h00f76863 /* 0x04b8 */;
            303: data_o = 32'h00813403 /* 0x04bc */;
            304: data_o = 32'h01010113 /* 0x04c0 */;
            305: data_o = 32'h00008067 /* 0x04c4 */;
            306: data_o = 32'hb0002773 /* 0x04c8 */;
            307: data_o = 32'hfedff06f /* 0x04cc */;
            308: data_o = 32'hf8010113 /* 0x04d0 */;
            309: data_o = 32'h06813823 /* 0x04d4 */;
            310: data_o = 32'h06113c23 /* 0x04d8 */;
            311: data_o = 32'h06913423 /* 0x04dc */;
            312: data_o = 32'h07213023 /* 0x04e0 */;
            313: data_o = 32'h05313c23 /* 0x04e4 */;
            314: data_o = 32'h05413823 /* 0x04e8 */;
            315: data_o = 32'h05513423 /* 0x04ec */;
            316: data_o = 32'h05613023 /* 0x04f0 */;
            317: data_o = 32'h03713c23 /* 0x04f4 */;
            318: data_o = 32'h03813823 /* 0x04f8 */;
            319: data_o = 32'h03913423 /* 0x04fc */;
            320: data_o = 32'h08010413 /* 0x0500 */;
            321: data_o = 32'hf15027f3 /* 0x0504 */;
            322: data_o = 32'hf8f42623 /* 0x0508 */;
            323: data_o = 32'h01002797 /* 0x050c */;
            324: data_o = 32'hae078c23 /* 0x0510 */;
            325: data_o = 32'hf8000793 /* 0x0514 */;
            326: data_o = 32'h01002717 /* 0x0518 */;
            327: data_o = 32'haef70a23 /* 0x051c */;
            328: data_o = 32'h00300793 /* 0x0520 */;
            329: data_o = 32'h01002717 /* 0x0524 */;
            330: data_o = 32'hacf70e23 /* 0x0528 */;
            331: data_o = 32'h01002717 /* 0x052c */;
            332: data_o = 32'hac070c23 /* 0x0530 */;
            333: data_o = 32'h01002717 /* 0x0534 */;
            334: data_o = 32'hacf70c23 /* 0x0538 */;
            335: data_o = 32'hfc700793 /* 0x053c */;
            336: data_o = 32'h01002717 /* 0x0540 */;
            337: data_o = 32'hacf70423 /* 0x0544 */;
            338: data_o = 32'h00100913 /* 0x0548 */;
            339: data_o = 32'h02200793 /* 0x054c */;
            340: data_o = 32'h01002717 /* 0x0550 */;
            341: data_o = 32'hacf70023 /* 0x0554 */;
            342: data_o = 32'h01f91993 /* 0x0558 */;
            343: data_o = 32'h00000a17 /* 0x055c */;
            344: data_o = 32'h28ca0a13 /* 0x0560 */;
            345: data_o = 32'h00000a97 /* 0x0564 */;
            346: data_o = 32'h28ca8a93 /* 0x0568 */;
            347: data_o = 32'h00000b17 /* 0x056c */;
            348: data_o = 32'h2a4b0b13 /* 0x0570 */;
            349: data_o = 32'h00000b97 /* 0x0574 */;
            350: data_o = 32'h2a4b8b93 /* 0x0578 */;
            351: data_o = 32'h000a0593 /* 0x057c */;
            352: data_o = 32'h00000513 /* 0x0580 */;
            353: data_o = 32'hf9343823 /* 0x0584 */;
            354: data_o = 32'hb81ff0ef /* 0x0588 */;
            355: data_o = 32'h000a8593 /* 0x058c */;
            356: data_o = 32'h00000513 /* 0x0590 */;
            357: data_o = 32'hb75ff0ef /* 0x0594 */;
            358: data_o = 32'h000b0593 /* 0x0598 */;
            359: data_o = 32'h00000513 /* 0x059c */;
            360: data_o = 32'hb69ff0ef /* 0x05a0 */;
            361: data_o = 32'h000b8593 /* 0x05a4 */;
            362: data_o = 32'h00000513 /* 0x05a8 */;
            363: data_o = 32'hb5dff0ef /* 0x05ac */;
            364: data_o = 32'h00000613 /* 0x05b0 */;
            365: data_o = 32'h00100593 /* 0x05b4 */;
            366: data_o = 32'hf8c40513 /* 0x05b8 */;
            367: data_o = 32'hbb5ff0ef /* 0x05bc */;
            368: data_o = 32'h00000597 /* 0x05c0 */;
            369: data_o = 32'h26858593 /* 0x05c4 */;
            370: data_o = 32'h00000513 /* 0x05c8 */;
            371: data_o = 32'hb3dff0ef /* 0x05cc */;
            372: data_o = 32'h00000597 /* 0x05d0 */;
            373: data_o = 32'h28858593 /* 0x05d4 */;
            374: data_o = 32'h00000513 /* 0x05d8 */;
            375: data_o = 32'hb2dff0ef /* 0x05dc */;
            376: data_o = 32'h00000597 /* 0x05e0 */;
            377: data_o = 32'h29058593 /* 0x05e4 */;
            378: data_o = 32'h00000513 /* 0x05e8 */;
            379: data_o = 32'hb1dff0ef /* 0x05ec */;
            380: data_o = 32'h00000613 /* 0x05f0 */;
            381: data_o = 32'h00800593 /* 0x05f4 */;
            382: data_o = 32'hf9040513 /* 0x05f8 */;
            383: data_o = 32'hb75ff0ef /* 0x05fc */;
            384: data_o = 32'h00000597 /* 0x0600 */;
            385: data_o = 32'h29058593 /* 0x0604 */;
            386: data_o = 32'h00000513 /* 0x0608 */;
            387: data_o = 32'hafdff0ef /* 0x060c */;
            388: data_o = 32'h00000613 /* 0x0610 */;
            389: data_o = 32'h00800593 /* 0x0614 */;
            390: data_o = 32'hf9040513 /* 0x0618 */;
            391: data_o = 32'hb55ff0ef /* 0x061c */;
            392: data_o = 32'h00000597 /* 0x0620 */;
            393: data_o = 32'h29058593 /* 0x0624 */;
            394: data_o = 32'h00000513 /* 0x0628 */;
            395: data_o = 32'haddff0ef /* 0x062c */;
            396: data_o = 32'h00000613 /* 0x0630 */;
            397: data_o = 32'h00800593 /* 0x0634 */;
            398: data_o = 32'hf9040513 /* 0x0638 */;
            399: data_o = 32'hb35ff0ef /* 0x063c */;
            400: data_o = 32'h00000513 /* 0x0640 */;
            401: data_o = 32'ha85ff0ef /* 0x0644 */;
            402: data_o = 32'hfcf5051b /* 0x0648 */;
            403: data_o = 32'h09250e63 /* 0x064c */;
            404: data_o = 32'h02a94263 /* 0x0650 */;
            405: data_o = 32'hf20514e3 /* 0x0654 */;
            406: data_o = 32'h00000597 /* 0x0658 */;
            407: data_o = 32'h27858593 /* 0x065c */;
            408: data_o = 32'h00000513 /* 0x0660 */;
            409: data_o = 32'haa5ff0ef /* 0x0664 */;
            410: data_o = 32'hf1402573 /* 0x0668 */;
            411: data_o = 32'h00100073 /* 0x066c */;
            412: data_o = 32'hf0dff06f /* 0x0670 */;
            413: data_o = 32'h00200793 /* 0x0674 */;
            414: data_o = 32'h08f50e63 /* 0x0678 */;
            415: data_o = 32'h00300793 /* 0x067c */;
            416: data_o = 32'heef51ee3 /* 0x0680 */;
            417: data_o = 32'h00000597 /* 0x0684 */;
            418: data_o = 32'h2dc58593 /* 0x0688 */;
            419: data_o = 32'h00000513 /* 0x068c */;
            420: data_o = 32'ha79ff0ef /* 0x0690 */;
            421: data_o = 32'hf9040513 /* 0x0694 */;
            422: data_o = 32'h00000613 /* 0x0698 */;
            423: data_o = 32'h00800593 /* 0x069c */;
            424: data_o = 32'had1ff0ef /* 0x06a0 */;
            425: data_o = 32'h00000597 /* 0x06a4 */;
            426: data_o = 32'h2d458593 /* 0x06a8 */;
            427: data_o = 32'h00000513 /* 0x06ac */;
            428: data_o = 32'ha59ff0ef /* 0x06b0 */;
            429: data_o = 32'h07813083 /* 0x06b4 */;
            430: data_o = 32'h07013403 /* 0x06b8 */;
            431: data_o = 32'h06813483 /* 0x06bc */;
            432: data_o = 32'h06013903 /* 0x06c0 */;
            433: data_o = 32'h05813983 /* 0x06c4 */;
            434: data_o = 32'h05013a03 /* 0x06c8 */;
            435: data_o = 32'h04813a83 /* 0x06cc */;
            436: data_o = 32'h04013b03 /* 0x06d0 */;
            437: data_o = 32'h03813b83 /* 0x06d4 */;
            438: data_o = 32'h03013c03 /* 0x06d8 */;
            439: data_o = 32'h02813c83 /* 0x06dc */;
            440: data_o = 32'h08010113 /* 0x06e0 */;
            441: data_o = 32'h00008067 /* 0x06e4 */;
            442: data_o = 32'h02faf537 /* 0x06e8 */;
            443: data_o = 32'h08050513 /* 0x06ec */;
            444: data_o = 32'hdb5ff0ef /* 0x06f0 */;
            445: data_o = 32'hf9043583 /* 0x06f4 */;
            446: data_o = 32'h00000513 /* 0x06f8 */;
            447: data_o = 32'hc4dff0ef /* 0x06fc */;
            448: data_o = 32'h00000597 /* 0x0700 */;
            449: data_o = 32'h0d058593 /* 0x0704 */;
            450: data_o = 32'h00000513 /* 0x0708 */;
            451: data_o = 32'h9fdff0ef /* 0x070c */;
            452: data_o = 32'he6dff06f /* 0x0710 */;
            453: data_o = 32'h00000597 /* 0x0714 */;
            454: data_o = 32'h1e458593 /* 0x0718 */;
            455: data_o = 32'h00000513 /* 0x071c */;
            456: data_o = 32'hf9840c13 /* 0x0720 */;
            457: data_o = 32'h9e5ff0ef /* 0x0724 */;
            458: data_o = 32'h000c0493 /* 0x0728 */;
            459: data_o = 32'h00d00c93 /* 0x072c */;
            460: data_o = 32'h00000513 /* 0x0730 */;
            461: data_o = 32'h995ff0ef /* 0x0734 */;
            462: data_o = 32'h00ac0023 /* 0x0738 */;
            463: data_o = 32'h07951c63 /* 0x073c */;
            464: data_o = 32'h00048793 /* 0x0740 */;
            465: data_o = 32'h000c0023 /* 0x0744 */;
            466: data_o = 32'h00000493 /* 0x0748 */;
            467: data_o = 32'h00a00693 /* 0x074c */;
            468: data_o = 32'h0007c703 /* 0x0750 */;
            469: data_o = 32'h06071463 /* 0x0754 */;
            470: data_o = 32'h00000597 /* 0x0758 */;
            471: data_o = 32'h1d058593 /* 0x075c */;
            472: data_o = 32'h00000513 /* 0x0760 */;
            473: data_o = 32'h9a5ff0ef /* 0x0764 */;
            474: data_o = 32'h00000613 /* 0x0768 */;
            475: data_o = 32'hf9040513 /* 0x076c */;
            476: data_o = 32'h00800593 /* 0x0770 */;
            477: data_o = 32'h9fdff0ef /* 0x0774 */;
            478: data_o = 32'h00000597 /* 0x0778 */;
            479: data_o = 32'h1c858593 /* 0x077c */;
            480: data_o = 32'h00000513 /* 0x0780 */;
            481: data_o = 32'h985ff0ef /* 0x0784 */;
            482: data_o = 32'hf9043503 /* 0x0788 */;
            483: data_o = 32'h00100613 /* 0x078c */;
            484: data_o = 32'h0004859b /* 0x0790 */;
            485: data_o = 32'h9ddff0ef /* 0x0794 */;
            486: data_o = 32'h00000597 /* 0x0798 */;
            487: data_o = 32'h1b058593 /* 0x079c */;
            488: data_o = 32'h00000513 /* 0x07a0 */;
            489: data_o = 32'h965ff0ef /* 0x07a4 */;
            490: data_o = 32'h00000513 /* 0x07a8 */;
            491: data_o = 32'h91dff0ef /* 0x07ac */;
            492: data_o = 32'hdcdff06f /* 0x07b0 */;
            493: data_o = 32'h001c0c13 /* 0x07b4 */;
            494: data_o = 32'hf79ff06f /* 0x07b8 */;
            495: data_o = 32'h02d484b3 /* 0x07bc */;
            496: data_o = 32'h00178793 /* 0x07c0 */;
            497: data_o = 32'hfd048493 /* 0x07c4 */;
            498: data_o = 32'h009704b3 /* 0x07c8 */;
            499: data_o = 32'hf85ff06f /* 0x07cc */;
            500: data_o = 32'h20090a0d /* 0x07d0 */;
            501: data_o = 32'h64616f4c /* 0x07d4 */;
            502: data_o = 32'h6e696620 /* 0x07d8 */;
            503: data_o = 32'h65687369 /* 0x07dc */;
            504: data_o = 32'h0d202e64 /* 0x07e0 */;
            505: data_o = 32'h000a0d0a /* 0x07e4 */;
            506: data_o = 32'h4a325b1b /* 0x07e8 */;
            507: data_o = 32'h00000000 /* 0x07ec */;
            508: data_o = 32'h09090a0d /* 0x07f0 */;
            509: data_o = 32'h6c655720 /* 0x07f4 */;
            510: data_o = 32'h656d6f63 /* 0x07f8 */;
            511: data_o = 32'h206f7420 /* 0x07fc */;
            512: data_o = 32'h414d6548 /* 0x0800 */;
            513: data_o = 32'h42204169 /* 0x0804 */;
            514: data_o = 32'h72746f6f /* 0x0808 */;
            515: data_o = 32'h00006d6f /* 0x080c */;
            516: data_o = 32'h00000a0d /* 0x0810 */;
            517: data_o = 32'h00000000 /* 0x0814 */;
            518: data_o = 32'h20090a0d /* 0x0818 */;
            519: data_o = 32'h70696843 /* 0x081c */;
            520: data_o = 32'h3a444920 /* 0x0820 */;
            521: data_o = 32'h00783020 /* 0x0824 */;
            522: data_o = 32'h20090a0d /* 0x0828 */;
            523: data_o = 32'h65746e45 /* 0x082c */;
            524: data_o = 32'h68742072 /* 0x0830 */;
            525: data_o = 32'h756e2065 /* 0x0834 */;
            526: data_o = 32'h7265626d /* 0x0838 */;
            527: data_o = 32'h206f7420 /* 0x083c */;
            528: data_o = 32'h656c6573 /* 0x0840 */;
            529: data_o = 32'h74207463 /* 0x0844 */;
            530: data_o = 32'h6d206568 /* 0x0848 */;
            531: data_o = 32'h3a65646f /* 0x084c */;
            532: data_o = 32'h00000020 /* 0x0850 */;
            533: data_o = 32'h00000000 /* 0x0854 */;
            534: data_o = 32'h20090a0d /* 0x0858 */;
            535: data_o = 32'h4c202e31 /* 0x085c */;
            536: data_o = 32'h2064616f /* 0x0860 */;
            537: data_o = 32'h6d6f7266 /* 0x0864 */;
            538: data_o = 32'h41544a20 /* 0x0868 */;
            539: data_o = 32'h00000047 /* 0x086c */;
            540: data_o = 32'h20090a0d /* 0x0870 */;
            541: data_o = 32'h4c202e32 /* 0x0874 */;
            542: data_o = 32'h2064616f /* 0x0878 */;
            543: data_o = 32'h6d6f7266 /* 0x087c */;
            544: data_o = 32'h52415520 /* 0x0880 */;
            545: data_o = 32'h6f742054 /* 0x0884 */;
            546: data_o = 32'h00783020 /* 0x0888 */;
            547: data_o = 32'h00000000 /* 0x088c */;
            548: data_o = 32'h20090a0d /* 0x0890 */;
            549: data_o = 32'h50202e33 /* 0x0894 */;
            550: data_o = 32'h746e6972 /* 0x0898 */;
            551: data_o = 32'h6d656d20 /* 0x089c */;
            552: data_o = 32'h2079726f /* 0x08a0 */;
            553: data_o = 32'h6d6f7266 /* 0x08a4 */;
            554: data_o = 32'h00783020 /* 0x08a8 */;
            555: data_o = 32'h00000000 /* 0x08ac */;
            556: data_o = 32'h20090a0d /* 0x08b0 */;
            557: data_o = 32'h43202e34 /* 0x08b4 */;
            558: data_o = 32'h69746e6f /* 0x08b8 */;
            559: data_o = 32'h2065756e /* 0x08bc */;
            560: data_o = 32'h42206f74 /* 0x08c0 */;
            561: data_o = 32'h20746f6f /* 0x08c4 */;
            562: data_o = 32'h6d6f7266 /* 0x08c8 */;
            563: data_o = 32'h00783020 /* 0x08cc */;
            564: data_o = 32'h20090a0d /* 0x08d0 */;
            565: data_o = 32'h646e6148 /* 0x08d4 */;
            566: data_o = 32'h7265766f /* 0x08d8 */;
            567: data_o = 32'h206f7420 /* 0x08dc */;
            568: data_o = 32'h75626564 /* 0x08e0 */;
            569: data_o = 32'h72656767 /* 0x08e4 */;
            570: data_o = 32'h202e2e2e /* 0x08e8 */;
            571: data_o = 32'h0a0d0a0d /* 0x08ec */;
            572: data_o = 32'h00000000 /* 0x08f0 */;
            573: data_o = 32'h00000000 /* 0x08f4 */;
            574: data_o = 32'h20090a0d /* 0x08f8 */;
            575: data_o = 32'h65746e45 /* 0x08fc */;
            576: data_o = 32'h68742072 /* 0x0900 */;
            577: data_o = 32'h69732065 /* 0x0904 */;
            578: data_o = 32'h6f20657a /* 0x0908 */;
            579: data_o = 32'h68742066 /* 0x090c */;
            580: data_o = 32'h656d2065 /* 0x0910 */;
            581: data_o = 32'h79726f6d /* 0x0914 */;
            582: data_o = 32'h206e6920 /* 0x0918 */;
            583: data_o = 32'h65747962 /* 0x091c */;
            584: data_o = 32'h0000203a /* 0x0920 */;
            585: data_o = 32'h00000000 /* 0x0924 */;
            586: data_o = 32'h20090a0d /* 0x0928 */;
            587: data_o = 32'h20656854 /* 0x092c */;
            588: data_o = 32'h6f6d656d /* 0x0930 */;
            589: data_o = 32'h66207972 /* 0x0934 */;
            590: data_o = 32'h206d6f72 /* 0x0938 */;
            591: data_o = 32'h00007830 /* 0x093c */;
            592: data_o = 32'h003a7369 /* 0x0940 */;
            593: data_o = 32'h00000000 /* 0x0944 */;
            594: data_o = 32'h0a0d0a0d /* 0x0948 */;
            595: data_o = 32'h72502009 /* 0x094c */;
            596: data_o = 32'h20746e69 /* 0x0950 */;
            597: data_o = 32'h696e6966 /* 0x0954 */;
            598: data_o = 32'h64656873 /* 0x0958 */;
            599: data_o = 32'h0000202e /* 0x095c */;
            600: data_o = 32'h20090a0d /* 0x0960 */;
            601: data_o = 32'h746f6f42 /* 0x0964 */;
            602: data_o = 32'h20676e69 /* 0x0968 */;
            603: data_o = 32'h30207461 /* 0x096c */;
            604: data_o = 32'h00000078 /* 0x0970 */;
            605: data_o = 32'h00000000 /* 0x0974 */;
            606: data_o = 32'h0d2e2e2e /* 0x0978 */;
            607: data_o = 32'h000a0d0a /* 0x097c */;
            608: data_o = 32'h33323130 /* 0x0980 */;
            609: data_o = 32'h37363534 /* 0x0984 */;
            610: data_o = 32'h42413938 /* 0x0988 */;
            611: data_o = 32'h46454443 /* 0x098c */;
            612: data_o = 32'h00000000 /* 0x0990 */;
            613: data_o = 32'h00000000 /* 0x0994 */;
            614: data_o = 32'h00000000 /* 0x0998 */;
            615: data_o = 32'h00000000 /* 0x099c */;
            616: data_o = 32'h00000000 /* 0x09a0 */;
            617: data_o = 32'h00000000 /* 0x09a4 */;
            618: data_o = 32'h00000000 /* 0x09a8 */;
            619: data_o = 32'h00000000 /* 0x09ac */;
            620: data_o = 32'h00000000 /* 0x09b0 */;
            621: data_o = 32'h00000000 /* 0x09b4 */;
            622: data_o = 32'h00000000 /* 0x09b8 */;
            623: data_o = 32'h00000000 /* 0x09bc */;
            624: data_o = 32'h00000000 /* 0x09c0 */;
            625: data_o = 32'h00000000 /* 0x09c4 */;
            626: data_o = 32'h00000000 /* 0x09c8 */;
            627: data_o = 32'h00000000 /* 0x09cc */;
            628: data_o = 32'h00000000 /* 0x09d0 */;
            629: data_o = 32'h00000000 /* 0x09d4 */;
            630: data_o = 32'h00000000 /* 0x09d8 */;
            631: data_o = 32'h00000000 /* 0x09dc */;
            632: data_o = 32'h00000000 /* 0x09e0 */;
            633: data_o = 32'h00000000 /* 0x09e4 */;
            634: data_o = 32'h00000000 /* 0x09e8 */;
            635: data_o = 32'h00000000 /* 0x09ec */;
            636: data_o = 32'h00000000 /* 0x09f0 */;
            637: data_o = 32'h00000000 /* 0x09f4 */;
            638: data_o = 32'h00000000 /* 0x09f8 */;
            639: data_o = 32'h00000000 /* 0x09fc */;
            640: data_o = 32'h00000000 /* 0x0a00 */;
            641: data_o = 32'h00000000 /* 0x0a04 */;
            642: data_o = 32'h00000000 /* 0x0a08 */;
            643: data_o = 32'h00000000 /* 0x0a0c */;
            644: data_o = 32'h00000000 /* 0x0a10 */;
            645: data_o = 32'h00000000 /* 0x0a14 */;
            646: data_o = 32'h00000000 /* 0x0a18 */;
            647: data_o = 32'h00000000 /* 0x0a1c */;
            648: data_o = 32'h00000000 /* 0x0a20 */;
            649: data_o = 32'h00000000 /* 0x0a24 */;
            650: data_o = 32'h00000000 /* 0x0a28 */;
            651: data_o = 32'h00000000 /* 0x0a2c */;
            652: data_o = 32'h00000000 /* 0x0a30 */;
            653: data_o = 32'h00000000 /* 0x0a34 */;
            654: data_o = 32'h00000000 /* 0x0a38 */;
            655: data_o = 32'h00000000 /* 0x0a3c */;
            656: data_o = 32'h00000000 /* 0x0a40 */;
            657: data_o = 32'h00000000 /* 0x0a44 */;
            658: data_o = 32'h00000000 /* 0x0a48 */;
            659: data_o = 32'h00000000 /* 0x0a4c */;
            660: data_o = 32'h00000000 /* 0x0a50 */;
            661: data_o = 32'h00000000 /* 0x0a54 */;
            662: data_o = 32'h00000000 /* 0x0a58 */;
            663: data_o = 32'h00000000 /* 0x0a5c */;
            664: data_o = 32'h00000000 /* 0x0a60 */;
            665: data_o = 32'h00000000 /* 0x0a64 */;
            666: data_o = 32'h00000000 /* 0x0a68 */;
            667: data_o = 32'h00000000 /* 0x0a6c */;
            668: data_o = 32'h00000000 /* 0x0a70 */;
            669: data_o = 32'h00000000 /* 0x0a74 */;
            670: data_o = 32'h00000000 /* 0x0a78 */;
            671: data_o = 32'h00000000 /* 0x0a7c */;
            672: data_o = 32'h00000000 /* 0x0a80 */;
            673: data_o = 32'h00000000 /* 0x0a84 */;
            674: data_o = 32'h00000000 /* 0x0a88 */;
            675: data_o = 32'h00000000 /* 0x0a8c */;
            676: data_o = 32'h00000000 /* 0x0a90 */;
            677: data_o = 32'h00000000 /* 0x0a94 */;
            678: data_o = 32'h00000000 /* 0x0a98 */;
            679: data_o = 32'h00000000 /* 0x0a9c */;
            680: data_o = 32'h00000000 /* 0x0aa0 */;
            681: data_o = 32'h00000000 /* 0x0aa4 */;
            682: data_o = 32'h00000000 /* 0x0aa8 */;
            683: data_o = 32'h00000000 /* 0x0aac */;
            684: data_o = 32'h00000000 /* 0x0ab0 */;
            685: data_o = 32'h00000000 /* 0x0ab4 */;
            686: data_o = 32'h00000000 /* 0x0ab8 */;
            687: data_o = 32'h00000000 /* 0x0abc */;
            688: data_o = 32'h00000000 /* 0x0ac0 */;
            689: data_o = 32'h00000000 /* 0x0ac4 */;
            690: data_o = 32'h00000000 /* 0x0ac8 */;
            691: data_o = 32'h00000000 /* 0x0acc */;
            692: data_o = 32'h00000000 /* 0x0ad0 */;
            693: data_o = 32'h00000000 /* 0x0ad4 */;
            694: data_o = 32'h00000000 /* 0x0ad8 */;
            695: data_o = 32'h00000000 /* 0x0adc */;
            696: data_o = 32'h00000000 /* 0x0ae0 */;
            697: data_o = 32'h00000000 /* 0x0ae4 */;
            698: data_o = 32'h00000000 /* 0x0ae8 */;
            699: data_o = 32'h00000000 /* 0x0aec */;
            700: data_o = 32'h00000000 /* 0x0af0 */;
            701: data_o = 32'h00000000 /* 0x0af4 */;
            702: data_o = 32'h00000000 /* 0x0af8 */;
            703: data_o = 32'h00000000 /* 0x0afc */;
            704: data_o = 32'h00000000 /* 0x0b00 */;
            705: data_o = 32'h00000000 /* 0x0b04 */;
            706: data_o = 32'h00000000 /* 0x0b08 */;
            707: data_o = 32'h00000000 /* 0x0b0c */;
            708: data_o = 32'h00000000 /* 0x0b10 */;
            709: data_o = 32'h00000000 /* 0x0b14 */;
            710: data_o = 32'h00000000 /* 0x0b18 */;
            711: data_o = 32'h00000000 /* 0x0b1c */;
            712: data_o = 32'h00000000 /* 0x0b20 */;
            713: data_o = 32'h00000000 /* 0x0b24 */;
            714: data_o = 32'h00000000 /* 0x0b28 */;
            715: data_o = 32'h00000000 /* 0x0b2c */;
            716: data_o = 32'h00000000 /* 0x0b30 */;
            717: data_o = 32'h00000000 /* 0x0b34 */;
            718: data_o = 32'h00000000 /* 0x0b38 */;
            719: data_o = 32'h00000000 /* 0x0b3c */;
            720: data_o = 32'h00000000 /* 0x0b40 */;
            721: data_o = 32'h00000000 /* 0x0b44 */;
            722: data_o = 32'h00000000 /* 0x0b48 */;
            723: data_o = 32'h00000000 /* 0x0b4c */;
            724: data_o = 32'h00000000 /* 0x0b50 */;
            725: data_o = 32'h00000000 /* 0x0b54 */;
            726: data_o = 32'h00000000 /* 0x0b58 */;
            727: data_o = 32'h00000000 /* 0x0b5c */;
            728: data_o = 32'h00000000 /* 0x0b60 */;
            729: data_o = 32'h00000000 /* 0x0b64 */;
            730: data_o = 32'h00000000 /* 0x0b68 */;
            731: data_o = 32'h00000000 /* 0x0b6c */;
            732: data_o = 32'h00000000 /* 0x0b70 */;
            733: data_o = 32'h00000000 /* 0x0b74 */;
            734: data_o = 32'h00000000 /* 0x0b78 */;
            735: data_o = 32'h00000000 /* 0x0b7c */;
            736: data_o = 32'h00000000 /* 0x0b80 */;
            737: data_o = 32'h00000000 /* 0x0b84 */;
            738: data_o = 32'h00000000 /* 0x0b88 */;
            739: data_o = 32'h00000000 /* 0x0b8c */;
            740: data_o = 32'h00000000 /* 0x0b90 */;
            741: data_o = 32'h00000000 /* 0x0b94 */;
            742: data_o = 32'h00000000 /* 0x0b98 */;
            743: data_o = 32'h00000000 /* 0x0b9c */;
            744: data_o = 32'h00000000 /* 0x0ba0 */;
            745: data_o = 32'h00000000 /* 0x0ba4 */;
            746: data_o = 32'h00000000 /* 0x0ba8 */;
            747: data_o = 32'h00000000 /* 0x0bac */;
            748: data_o = 32'h00000000 /* 0x0bb0 */;
            749: data_o = 32'h00000000 /* 0x0bb4 */;
            750: data_o = 32'h00000000 /* 0x0bb8 */;
            751: data_o = 32'h00000000 /* 0x0bbc */;
            752: data_o = 32'h00000000 /* 0x0bc0 */;
            753: data_o = 32'h00000000 /* 0x0bc4 */;
            754: data_o = 32'h00000000 /* 0x0bc8 */;
            755: data_o = 32'h00000000 /* 0x0bcc */;
            756: data_o = 32'h00000000 /* 0x0bd0 */;
            757: data_o = 32'h00000000 /* 0x0bd4 */;
            758: data_o = 32'h00000000 /* 0x0bd8 */;
            759: data_o = 32'h00000000 /* 0x0bdc */;
            760: data_o = 32'h00000000 /* 0x0be0 */;
            761: data_o = 32'h00000000 /* 0x0be4 */;
            762: data_o = 32'h00000000 /* 0x0be8 */;
            763: data_o = 32'h00000000 /* 0x0bec */;
            764: data_o = 32'h00000000 /* 0x0bf0 */;
            765: data_o = 32'h00000000 /* 0x0bf4 */;
            766: data_o = 32'h00000000 /* 0x0bf8 */;
            767: data_o = 32'h00000000 /* 0x0bfc */;
            768: data_o = 32'h00000000 /* 0x0c00 */;
            769: data_o = 32'h00000000 /* 0x0c04 */;
            770: data_o = 32'h00000000 /* 0x0c08 */;
            771: data_o = 32'h00000000 /* 0x0c0c */;
            772: data_o = 32'h00000000 /* 0x0c10 */;
            773: data_o = 32'h00000000 /* 0x0c14 */;
            774: data_o = 32'h00000000 /* 0x0c18 */;
            775: data_o = 32'h00000000 /* 0x0c1c */;
            776: data_o = 32'h00000000 /* 0x0c20 */;
            777: data_o = 32'h00000000 /* 0x0c24 */;
            778: data_o = 32'h00000000 /* 0x0c28 */;
            779: data_o = 32'h00000000 /* 0x0c2c */;
            780: data_o = 32'h00000000 /* 0x0c30 */;
            781: data_o = 32'h00000000 /* 0x0c34 */;
            782: data_o = 32'h00000000 /* 0x0c38 */;
            783: data_o = 32'h00000000 /* 0x0c3c */;
            784: data_o = 32'h00000000 /* 0x0c40 */;
            785: data_o = 32'h00000000 /* 0x0c44 */;
            786: data_o = 32'h00000000 /* 0x0c48 */;
            787: data_o = 32'h00000000 /* 0x0c4c */;
            788: data_o = 32'h00000000 /* 0x0c50 */;
            789: data_o = 32'h00000000 /* 0x0c54 */;
            790: data_o = 32'h00000000 /* 0x0c58 */;
            791: data_o = 32'h00000000 /* 0x0c5c */;
            792: data_o = 32'h00000000 /* 0x0c60 */;
            793: data_o = 32'h00000000 /* 0x0c64 */;
            794: data_o = 32'h00000000 /* 0x0c68 */;
            795: data_o = 32'h00000000 /* 0x0c6c */;
            796: data_o = 32'h00000000 /* 0x0c70 */;
            797: data_o = 32'h00000000 /* 0x0c74 */;
            798: data_o = 32'h00000000 /* 0x0c78 */;
            799: data_o = 32'h00000000 /* 0x0c7c */;
            800: data_o = 32'h00000000 /* 0x0c80 */;
            801: data_o = 32'h00000000 /* 0x0c84 */;
            802: data_o = 32'h00000000 /* 0x0c88 */;
            803: data_o = 32'h00000000 /* 0x0c8c */;
            804: data_o = 32'h00000000 /* 0x0c90 */;
            805: data_o = 32'h00000000 /* 0x0c94 */;
            806: data_o = 32'h00000000 /* 0x0c98 */;
            807: data_o = 32'h00000000 /* 0x0c9c */;
            808: data_o = 32'h00000000 /* 0x0ca0 */;
            809: data_o = 32'h00000000 /* 0x0ca4 */;
            810: data_o = 32'h00000000 /* 0x0ca8 */;
            811: data_o = 32'h00000000 /* 0x0cac */;
            812: data_o = 32'h00000000 /* 0x0cb0 */;
            813: data_o = 32'h00000000 /* 0x0cb4 */;
            814: data_o = 32'h00000000 /* 0x0cb8 */;
            815: data_o = 32'h00000000 /* 0x0cbc */;
            816: data_o = 32'h00000000 /* 0x0cc0 */;
            817: data_o = 32'h00000000 /* 0x0cc4 */;
            818: data_o = 32'h00000000 /* 0x0cc8 */;
            819: data_o = 32'h00000000 /* 0x0ccc */;
            820: data_o = 32'h00000000 /* 0x0cd0 */;
            821: data_o = 32'h00000000 /* 0x0cd4 */;
            822: data_o = 32'h00000000 /* 0x0cd8 */;
            823: data_o = 32'h00000000 /* 0x0cdc */;
            824: data_o = 32'h00000000 /* 0x0ce0 */;
            825: data_o = 32'h00000000 /* 0x0ce4 */;
            826: data_o = 32'h00000000 /* 0x0ce8 */;
            827: data_o = 32'h00000000 /* 0x0cec */;
            828: data_o = 32'h00000000 /* 0x0cf0 */;
            829: data_o = 32'h00000000 /* 0x0cf4 */;
            830: data_o = 32'h00000000 /* 0x0cf8 */;
            831: data_o = 32'h00000000 /* 0x0cfc */;
            832: data_o = 32'h00000000 /* 0x0d00 */;
            833: data_o = 32'h00000000 /* 0x0d04 */;
            834: data_o = 32'h00000000 /* 0x0d08 */;
            835: data_o = 32'h00000000 /* 0x0d0c */;
            836: data_o = 32'h00000000 /* 0x0d10 */;
            837: data_o = 32'h00000000 /* 0x0d14 */;
            838: data_o = 32'h00000000 /* 0x0d18 */;
            839: data_o = 32'h00000000 /* 0x0d1c */;
            840: data_o = 32'h00000000 /* 0x0d20 */;
            841: data_o = 32'h00000000 /* 0x0d24 */;
            842: data_o = 32'h00000000 /* 0x0d28 */;
            843: data_o = 32'h00000000 /* 0x0d2c */;
            844: data_o = 32'h00000000 /* 0x0d30 */;
            845: data_o = 32'h00000000 /* 0x0d34 */;
            846: data_o = 32'h00000000 /* 0x0d38 */;
            847: data_o = 32'h00000000 /* 0x0d3c */;
            848: data_o = 32'h00000000 /* 0x0d40 */;
            849: data_o = 32'h00000000 /* 0x0d44 */;
            850: data_o = 32'h00000000 /* 0x0d48 */;
            851: data_o = 32'h00000000 /* 0x0d4c */;
            852: data_o = 32'h00000000 /* 0x0d50 */;
            853: data_o = 32'h00000000 /* 0x0d54 */;
            854: data_o = 32'h00000000 /* 0x0d58 */;
            855: data_o = 32'h00000000 /* 0x0d5c */;
            856: data_o = 32'h00000000 /* 0x0d60 */;
            857: data_o = 32'h00000000 /* 0x0d64 */;
            858: data_o = 32'h00000000 /* 0x0d68 */;
            859: data_o = 32'h00000000 /* 0x0d6c */;
            860: data_o = 32'h00000000 /* 0x0d70 */;
            861: data_o = 32'h00000000 /* 0x0d74 */;
            862: data_o = 32'h00000000 /* 0x0d78 */;
            863: data_o = 32'h00000000 /* 0x0d7c */;
            864: data_o = 32'h00000000 /* 0x0d80 */;
            865: data_o = 32'h00000000 /* 0x0d84 */;
            866: data_o = 32'h00000000 /* 0x0d88 */;
            867: data_o = 32'h00000000 /* 0x0d8c */;
            868: data_o = 32'h00000000 /* 0x0d90 */;
            869: data_o = 32'h00000000 /* 0x0d94 */;
            870: data_o = 32'h00000000 /* 0x0d98 */;
            871: data_o = 32'h00000000 /* 0x0d9c */;
            872: data_o = 32'h00000000 /* 0x0da0 */;
            873: data_o = 32'h00000000 /* 0x0da4 */;
            874: data_o = 32'h00000000 /* 0x0da8 */;
            875: data_o = 32'h00000000 /* 0x0dac */;
            876: data_o = 32'h00000000 /* 0x0db0 */;
            877: data_o = 32'h00000000 /* 0x0db4 */;
            878: data_o = 32'h00000000 /* 0x0db8 */;
            879: data_o = 32'h00000000 /* 0x0dbc */;
            880: data_o = 32'h00000000 /* 0x0dc0 */;
            881: data_o = 32'h00000000 /* 0x0dc4 */;
            882: data_o = 32'h00000000 /* 0x0dc8 */;
            883: data_o = 32'h00000000 /* 0x0dcc */;
            884: data_o = 32'h00000000 /* 0x0dd0 */;
            885: data_o = 32'h00000000 /* 0x0dd4 */;
            886: data_o = 32'h00000000 /* 0x0dd8 */;
            887: data_o = 32'h00000000 /* 0x0ddc */;
            888: data_o = 32'h00000000 /* 0x0de0 */;
            889: data_o = 32'h00000000 /* 0x0de4 */;
            890: data_o = 32'h00000000 /* 0x0de8 */;
            891: data_o = 32'h00000000 /* 0x0dec */;
            892: data_o = 32'h00000000 /* 0x0df0 */;
            893: data_o = 32'h00000000 /* 0x0df4 */;
            894: data_o = 32'h00000000 /* 0x0df8 */;
            895: data_o = 32'h00000000 /* 0x0dfc */;
            896: data_o = 32'h00000000 /* 0x0e00 */;
            897: data_o = 32'h00000000 /* 0x0e04 */;
            898: data_o = 32'h00000000 /* 0x0e08 */;
            899: data_o = 32'h00000000 /* 0x0e0c */;
            900: data_o = 32'h00000000 /* 0x0e10 */;
            901: data_o = 32'h00000000 /* 0x0e14 */;
            902: data_o = 32'h00000000 /* 0x0e18 */;
            903: data_o = 32'h00000000 /* 0x0e1c */;
            904: data_o = 32'h00000000 /* 0x0e20 */;
            905: data_o = 32'h00000000 /* 0x0e24 */;
            906: data_o = 32'h00000000 /* 0x0e28 */;
            907: data_o = 32'h00000000 /* 0x0e2c */;
            908: data_o = 32'h00000000 /* 0x0e30 */;
            909: data_o = 32'h00000000 /* 0x0e34 */;
            910: data_o = 32'h00000000 /* 0x0e38 */;
            911: data_o = 32'h00000000 /* 0x0e3c */;
            912: data_o = 32'h00000000 /* 0x0e40 */;
            913: data_o = 32'h00000000 /* 0x0e44 */;
            914: data_o = 32'h00000000 /* 0x0e48 */;
            915: data_o = 32'h00000000 /* 0x0e4c */;
            916: data_o = 32'h00000000 /* 0x0e50 */;
            917: data_o = 32'h00000000 /* 0x0e54 */;
            918: data_o = 32'h00000000 /* 0x0e58 */;
            919: data_o = 32'h00000000 /* 0x0e5c */;
            920: data_o = 32'h00000000 /* 0x0e60 */;
            921: data_o = 32'h00000000 /* 0x0e64 */;
            922: data_o = 32'h00000000 /* 0x0e68 */;
            923: data_o = 32'h00000000 /* 0x0e6c */;
            924: data_o = 32'h00000000 /* 0x0e70 */;
            925: data_o = 32'h00000000 /* 0x0e74 */;
            926: data_o = 32'h00000000 /* 0x0e78 */;
            927: data_o = 32'h00000000 /* 0x0e7c */;
            928: data_o = 32'h00000000 /* 0x0e80 */;
            929: data_o = 32'h00000000 /* 0x0e84 */;
            930: data_o = 32'h00000000 /* 0x0e88 */;
            931: data_o = 32'h00000000 /* 0x0e8c */;
            932: data_o = 32'h00000000 /* 0x0e90 */;
            933: data_o = 32'h00000000 /* 0x0e94 */;
            934: data_o = 32'h00000000 /* 0x0e98 */;
            935: data_o = 32'h00000000 /* 0x0e9c */;
            936: data_o = 32'h00000000 /* 0x0ea0 */;
            937: data_o = 32'h00000000 /* 0x0ea4 */;
            938: data_o = 32'h00000000 /* 0x0ea8 */;
            939: data_o = 32'h00000000 /* 0x0eac */;
            940: data_o = 32'h00000000 /* 0x0eb0 */;
            941: data_o = 32'h00000000 /* 0x0eb4 */;
            942: data_o = 32'h00000000 /* 0x0eb8 */;
            943: data_o = 32'h00000000 /* 0x0ebc */;
            944: data_o = 32'h00000000 /* 0x0ec0 */;
            945: data_o = 32'h00000000 /* 0x0ec4 */;
            946: data_o = 32'h00000000 /* 0x0ec8 */;
            947: data_o = 32'h00000000 /* 0x0ecc */;
            948: data_o = 32'h00000000 /* 0x0ed0 */;
            949: data_o = 32'h00000000 /* 0x0ed4 */;
            950: data_o = 32'h00000000 /* 0x0ed8 */;
            951: data_o = 32'h00000000 /* 0x0edc */;
            952: data_o = 32'h00000000 /* 0x0ee0 */;
            953: data_o = 32'h00000000 /* 0x0ee4 */;
            954: data_o = 32'h00000000 /* 0x0ee8 */;
            955: data_o = 32'h00000000 /* 0x0eec */;
            956: data_o = 32'h00000000 /* 0x0ef0 */;
            957: data_o = 32'h00000000 /* 0x0ef4 */;
            958: data_o = 32'h00000000 /* 0x0ef8 */;
            959: data_o = 32'h00000000 /* 0x0efc */;
            960: data_o = 32'h00000000 /* 0x0f00 */;
            961: data_o = 32'h00000000 /* 0x0f04 */;
            962: data_o = 32'h00000000 /* 0x0f08 */;
            963: data_o = 32'h00000000 /* 0x0f0c */;
            964: data_o = 32'h00000000 /* 0x0f10 */;
            965: data_o = 32'h00000000 /* 0x0f14 */;
            966: data_o = 32'h00000000 /* 0x0f18 */;
            967: data_o = 32'h00000000 /* 0x0f1c */;
            968: data_o = 32'h00000000 /* 0x0f20 */;
            969: data_o = 32'h00000000 /* 0x0f24 */;
            970: data_o = 32'h00000000 /* 0x0f28 */;
            971: data_o = 32'h00000000 /* 0x0f2c */;
            972: data_o = 32'h00000000 /* 0x0f30 */;
            973: data_o = 32'h00000000 /* 0x0f34 */;
            974: data_o = 32'h00000000 /* 0x0f38 */;
            975: data_o = 32'h00000000 /* 0x0f3c */;
            976: data_o = 32'h00000000 /* 0x0f40 */;
            977: data_o = 32'h00000000 /* 0x0f44 */;
            978: data_o = 32'h00000000 /* 0x0f48 */;
            979: data_o = 32'h00000000 /* 0x0f4c */;
            980: data_o = 32'h00000000 /* 0x0f50 */;
            981: data_o = 32'h00000000 /* 0x0f54 */;
            982: data_o = 32'h00000000 /* 0x0f58 */;
            983: data_o = 32'h00000000 /* 0x0f5c */;
            984: data_o = 32'h00000000 /* 0x0f60 */;
            985: data_o = 32'h00000000 /* 0x0f64 */;
            986: data_o = 32'h00000000 /* 0x0f68 */;
            987: data_o = 32'h00000000 /* 0x0f6c */;
            988: data_o = 32'h00000000 /* 0x0f70 */;
            989: data_o = 32'h00000000 /* 0x0f74 */;
            990: data_o = 32'h00000000 /* 0x0f78 */;
            991: data_o = 32'h00000000 /* 0x0f7c */;
            992: data_o = 32'h00000000 /* 0x0f80 */;
            993: data_o = 32'h00000000 /* 0x0f84 */;
            994: data_o = 32'h00000000 /* 0x0f88 */;
            995: data_o = 32'h00000000 /* 0x0f8c */;
            996: data_o = 32'h00000000 /* 0x0f90 */;
            997: data_o = 32'h00000000 /* 0x0f94 */;
            998: data_o = 32'h00000000 /* 0x0f98 */;
            999: data_o = 32'h00000000 /* 0x0f9c */;
            1000: data_o = 32'h00000000 /* 0x0fa0 */;
            1001: data_o = 32'h00000000 /* 0x0fa4 */;
            1002: data_o = 32'h00000000 /* 0x0fa8 */;
            1003: data_o = 32'h00000000 /* 0x0fac */;
            1004: data_o = 32'h00000000 /* 0x0fb0 */;
            1005: data_o = 32'h00000000 /* 0x0fb4 */;
            1006: data_o = 32'h00000000 /* 0x0fb8 */;
            1007: data_o = 32'h00000000 /* 0x0fbc */;
            1008: data_o = 32'h00000000 /* 0x0fc0 */;
            1009: data_o = 32'h00000000 /* 0x0fc4 */;
            1010: data_o = 32'h00000000 /* 0x0fc8 */;
            1011: data_o = 32'h00000000 /* 0x0fcc */;
            1012: data_o = 32'h00000000 /* 0x0fd0 */;
            1013: data_o = 32'h00000000 /* 0x0fd4 */;
            1014: data_o = 32'h00000000 /* 0x0fd8 */;
            1015: data_o = 32'h00000000 /* 0x0fdc */;
            1016: data_o = 32'h00000000 /* 0x0fe0 */;
            1017: data_o = 32'h00000000 /* 0x0fe4 */;
            1018: data_o = 32'h00000000 /* 0x0fe8 */;
            1019: data_o = 32'h00000000 /* 0x0fec */;
            1020: data_o = 32'h00000000 /* 0x0ff0 */;
            1021: data_o = 32'h00000000 /* 0x0ff4 */;
            1022: data_o = 32'h00000000 /* 0x0ff8 */;
            1023: data_o = 32'h00000000 /* 0x0ffc */;
            default: data_o = '0;
        endcase
    end

endmodule
