// Copyright 2026 KU Leuven.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51
// Yunhao Deng <yunhao.deng@kuleuven.be>

module hemaia_io_pad (
    inout wire CRBL_X1_Y4,
    inout wire CRBL_X1_Y3,
    inout wire CRBL_X2_Y3,
    inout wire CRBL_X2_Y2,
    inout wire CRBL_X1_Y2,
    inout wire CRBL_X3_Y3,
    inout wire CRBL_X4_Y4,
    inout wire CRBL_X1_Y1,
    inout wire CRBL_X2_Y4,
    inout wire CRBL_X4_Y2,
    inout wire CRBL_X5_Y2,
    inout wire CRBL_X2_Y1,
    inout wire CRBL_X3_Y1,
    inout wire CRBL_X3_Y2,
    inout wire CRBL_X4_Y1,
    inout wire CRBL_X5_Y1,
    inout wire CRBL_X0_Y0,
    inout wire CRBL_X0_Y4,
    inout wire CRBL_X0_Y1,
    inout wire CRBL_X0_Y3,
    inout wire CRBL_X3_Y0,
    inout wire CRBL_X2_Y0,
    inout wire CRBL_X1_Y0,
    inout wire CRBL_X5_Y0,
    inout wire CRBL_X4_Y0,
    inout wire CRBL_X0_Y2,
    inout wire CRBL_X3_Y4,
    inout wire CRBL_X4_Y3,
    inout wire CRBL_X5_Y4,
    inout wire CRBL_X5_Y3,
    inout wire CRBR_X3_Y2,
    inout wire CRBR_X3_Y3,
    inout wire CRBR_X3_Y4,
    inout wire CRBR_X3_Y5,
    inout wire CRBR_X2_Y3,
    inout wire CRBR_X1_Y4,
    inout wire CRBR_X0_Y3,
    inout wire CRBR_X2_Y5,
    inout wire CRBR_X2_Y4,
    inout wire CRBR_X0_Y2,
    inout wire CRBR_X2_Y1,
    inout wire CRBR_X1_Y2,
    inout wire CRBR_X1_Y1,
    inout wire CRBR_X2_Y2,
    inout wire CRBR_X0_Y1,
    inout wire CRBR_X3_Y1,
    inout wire CRBR_X1_Y5,
    inout wire CRBR_X4_Y0,
    inout wire CRBR_X0_Y0,
    inout wire CRBR_X3_Y0,
    inout wire CRBR_X1_Y0,
    inout wire CRBR_X4_Y3,
    inout wire CRBR_X4_Y2,
    inout wire CRBR_X4_Y1,
    inout wire CRBR_X4_Y5,
    inout wire CRBR_X4_Y4,
    inout wire CRBR_X2_Y0,
    inout wire CRBR_X0_Y5,
    inout wire CRBR_X0_Y4,
    inout wire CRBR_X1_Y3,
    inout wire CRTL_X4_Y4,
    inout wire CRTL_X3_Y4,
    inout wire CRTL_X2_Y0,
    inout wire CRTL_X2_Y1,
    inout wire CRTL_X1_Y4,
    inout wire CRTL_X1_Y3,
    inout wire CRTL_X1_Y1,
    inout wire CRTL_X1_Y2,
    inout wire CRTL_X1_Y0,
    inout wire CRTL_X2_Y4,
    inout wire CRTL_X2_Y3,
    inout wire CRTL_X2_Y2,
    inout wire CRTL_X3_Y3,
    inout wire CRTL_X4_Y3,
    inout wire CRTL_X3_Y2,
    inout wire CRTL_X4_Y2,
    inout wire CRTL_X4_Y1,
    inout wire CRTL_X3_Y1,
    inout wire CRTL_X4_Y5,
    inout wire CRTL_X3_Y5,
    inout wire CRTL_X2_Y5,
    inout wire CRTL_X1_Y5,
    inout wire CRTL_X0_Y5,
    inout wire CRTL_X0_Y4,
    inout wire CRTL_X0_Y3,
    inout wire CRTL_X0_Y2,
    inout wire CRTL_X0_Y1,
    inout wire CRTL_X0_Y0,
    inout wire CRTL_X3_Y0,
    inout wire CRTL_X4_Y0,
    inout wire CRTR_X2_Y3,
    inout wire CRTR_X1_Y3,
    inout wire CRTR_X0_Y3,
    inout wire CRTR_X1_Y2,
    inout wire CRTR_X2_Y2,
    inout wire CRTR_X3_Y2,
    inout wire CRTR_X0_Y1,
    inout wire CRTR_X1_Y1,
    inout wire CRTR_X3_Y0,
    inout wire CRTR_X3_Y1,
    inout wire CRTR_X0_Y2,
    inout wire CRTR_X4_Y0,
    inout wire CRTR_X4_Y1,
    inout wire CRTR_X4_Y2,
    inout wire CRTR_X4_Y3,
    inout wire CRTR_X3_Y3,
    inout wire CRTR_X5_Y4,
    inout wire CRTR_X4_Y4,
    inout wire CRTR_X3_Y4,
    inout wire CRTR_X2_Y4,
    inout wire CRTR_X1_Y4,
    inout wire CRTR_X0_Y4,
    inout wire CRTR_X5_Y3,
    inout wire CRTR_X5_Y2,
    inout wire CRTR_X5_Y1,
    inout wire CRTR_X5_Y0,
    inout wire CRTR_X2_Y1,
    inout wire CRTR_X0_Y0,
    inout wire CRTR_X1_Y0,
    inout wire CRTR_X2_Y0,
    inout wire M_X0_Y9,
    inout wire M_X8_Y9,
    inout wire M_X9_Y9,
    inout wire M_X1_Y9,
    inout wire M_X3_Y9,
    inout wire M_X2_Y9,
    inout wire M_X4_Y9,
    inout wire M_X6_Y9,
    inout wire M_X7_Y9,
    inout wire M_X5_Y9,
    inout wire M_X9_Y8,
    inout wire M_X9_Y7,
    inout wire M_X9_Y6,
    inout wire M_X9_Y5,
    inout wire M_X9_Y4,
    inout wire M_X9_Y3,
    inout wire M_X9_Y2,
    inout wire M_X9_Y1,
    inout wire M_X9_Y0,
    inout wire M_X0_Y8,
    inout wire M_X0_Y7,
    inout wire M_X0_Y6,
    inout wire M_X0_Y5,
    inout wire M_X0_Y4,
    inout wire M_X0_Y3,
    inout wire M_X0_Y2,
    inout wire M_X0_Y1,
    inout wire M_X0_Y0,
    inout wire M_X8_Y0,
    inout wire M_X1_Y0,
    inout wire M_X3_Y0,
    inout wire M_X2_Y0,
    inout wire M_X4_Y0,
    inout wire M_X6_Y0,
    inout wire M_X7_Y0,
    inout wire M_X5_Y0,
    inout wire D2DE_X5_Y6,
    inout wire D2DE_X5_Y7,
    inout wire D2DE_X5_Y8,
    inout wire D2DE_X5_Y9,
    inout wire D2DE_X5_Y10,
    inout wire D2DE_X5_Y1,
    inout wire D2DE_X5_Y2,
    inout wire D2DE_X5_Y3,
    inout wire D2DE_X5_Y4,
    inout wire D2DE_X5_Y5,
    inout wire D2DE_X5_Y0,
    inout wire D2DE_X4_Y8,
    inout wire D2DE_X4_Y7,
    inout wire D2DE_X4_Y6,
    inout wire D2DE_X3_Y6,
    inout wire D2DE_X2_Y6,
    inout wire D2DE_X1_Y6,
    inout wire D2DE_X0_Y6,
    inout wire D2DE_X4_Y5,
    inout wire D2DE_X3_Y5,
    inout wire D2DE_X2_Y5,
    inout wire D2DE_X1_Y5,
    inout wire D2DE_X4_Y4,
    inout wire D2DE_X3_Y4,
    inout wire D2DE_X2_Y4,
    inout wire D2DE_X1_Y4,
    inout wire D2DE_X4_Y3,
    inout wire D2DE_X4_Y2,
    inout wire D2DE_X4_Y1,
    inout wire D2DE_X0_Y4,
    inout wire D2DE_X0_Y5,
    inout wire D2DE_X4_Y0,
    inout wire D2DE_X0_Y0,
    inout wire D2DE_X0_Y1,
    inout wire D2DE_X0_Y2,
    inout wire D2DE_X0_Y3,
    inout wire D2DE_X1_Y0,
    inout wire D2DE_X1_Y1,
    inout wire D2DE_X1_Y2,
    inout wire D2DE_X1_Y3,
    inout wire D2DE_X2_Y0,
    inout wire D2DE_X2_Y1,
    inout wire D2DE_X2_Y2,
    inout wire D2DE_X2_Y3,
    inout wire D2DE_X3_Y0,
    inout wire D2DE_X3_Y1,
    inout wire D2DE_X3_Y2,
    inout wire D2DE_X3_Y3,
    inout wire D2DE_X0_Y7,
    inout wire D2DE_X0_Y8,
    inout wire D2DE_X0_Y9,
    inout wire D2DE_X0_Y10,
    inout wire D2DE_X1_Y7,
    inout wire D2DE_X1_Y8,
    inout wire D2DE_X1_Y9,
    inout wire D2DE_X1_Y10,
    inout wire D2DE_X2_Y7,
    inout wire D2DE_X2_Y8,
    inout wire D2DE_X2_Y9,
    inout wire D2DE_X2_Y10,
    inout wire D2DE_X3_Y7,
    inout wire D2DE_X3_Y8,
    inout wire D2DE_X3_Y9,
    inout wire D2DE_X3_Y10,
    inout wire D2DE_X4_Y10,
    inout wire D2DE_X4_Y9,
    inout wire D2DN_X0_Y5,
    inout wire D2DN_X1_Y5,
    inout wire D2DN_X2_Y5,
    inout wire D2DN_X0_Y0,
    inout wire D2DN_X1_Y0,
    inout wire D2DN_X7_Y1,
    inout wire D2DN_X7_Y2,
    inout wire D2DN_X7_Y3,
    inout wire D2DN_X7_Y4,
    inout wire D2DN_X8_Y1,
    inout wire D2DN_X8_Y2,
    inout wire D2DN_X8_Y3,
    inout wire D2DN_X8_Y4,
    inout wire D2DN_X9_Y1,
    inout wire D2DN_X9_Y2,
    inout wire D2DN_X9_Y3,
    inout wire D2DN_X9_Y4,
    inout wire D2DN_X10_Y1,
    inout wire D2DN_X10_Y2,
    inout wire D2DN_X10_Y3,
    inout wire D2DN_X10_Y4,
    inout wire D2DN_X0_Y1,
    inout wire D2DN_X0_Y2,
    inout wire D2DN_X0_Y3,
    inout wire D2DN_X0_Y4,
    inout wire D2DN_X1_Y1,
    inout wire D2DN_X1_Y2,
    inout wire D2DN_X1_Y3,
    inout wire D2DN_X1_Y4,
    inout wire D2DN_X2_Y1,
    inout wire D2DN_X2_Y2,
    inout wire D2DN_X2_Y3,
    inout wire D2DN_X2_Y4,
    inout wire D2DN_X3_Y1,
    inout wire D2DN_X3_Y2,
    inout wire D2DN_X3_Y3,
    inout wire D2DN_X3_Y4,
    inout wire D2DN_X9_Y5,
    inout wire D2DN_X10_Y5,
    inout wire D2DN_X9_Y0,
    inout wire D2DN_X10_Y0,
    inout wire D2DN_X2_Y0,
    inout wire D2DN_X4_Y0,
    inout wire D2DN_X4_Y1,
    inout wire D2DN_X4_Y2,
    inout wire D2DN_X3_Y0,
    inout wire D2DN_X5_Y0,
    inout wire D2DN_X5_Y3,
    inout wire D2DN_X5_Y4,
    inout wire D2DN_X7_Y0,
    inout wire D2DN_X6_Y1,
    inout wire D2DN_X5_Y1,
    inout wire D2DN_X6_Y3,
    inout wire D2DN_X8_Y0,
    inout wire D2DN_X6_Y0,
    inout wire D2DN_X6_Y2,
    inout wire D2DN_X6_Y4,
    inout wire D2DN_X5_Y5,
    inout wire D2DN_X6_Y5,
    inout wire D2DN_X4_Y3,
    inout wire D2DN_X4_Y4,
    inout wire D2DN_X8_Y5,
    inout wire D2DN_X7_Y5,
    inout wire D2DN_X4_Y5,
    inout wire D2DN_X3_Y5,
    inout wire D2DN_X5_Y2,
    inout wire D2DS_X0_Y0,
    inout wire D2DS_X1_Y0,
    inout wire D2DS_X8_Y0,
    inout wire D2DS_X9_Y0,
    inout wire D2DS_X4_Y0,
    inout wire D2DS_X5_Y0,
    inout wire D2DS_X7_Y0,
    inout wire D2DS_X6_Y0,
    inout wire D2DS_X3_Y0,
    inout wire D2DS_X2_Y0,
    inout wire D2DS_X10_Y0,
    inout wire D2DS_X0_Y1,
    inout wire D2DS_X1_Y1,
    inout wire D2DS_X7_Y2,
    inout wire D2DS_X7_Y3,
    inout wire D2DS_X7_Y4,
    inout wire D2DS_X7_Y5,
    inout wire D2DS_X8_Y2,
    inout wire D2DS_X8_Y3,
    inout wire D2DS_X8_Y4,
    inout wire D2DS_X8_Y5,
    inout wire D2DS_X9_Y2,
    inout wire D2DS_X9_Y3,
    inout wire D2DS_X9_Y4,
    inout wire D2DS_X9_Y5,
    inout wire D2DS_X10_Y2,
    inout wire D2DS_X10_Y3,
    inout wire D2DS_X10_Y4,
    inout wire D2DS_X10_Y5,
    inout wire D2DS_X0_Y2,
    inout wire D2DS_X0_Y3,
    inout wire D2DS_X0_Y4,
    inout wire D2DS_X0_Y5,
    inout wire D2DS_X1_Y2,
    inout wire D2DS_X1_Y3,
    inout wire D2DS_X1_Y4,
    inout wire D2DS_X1_Y5,
    inout wire D2DS_X2_Y2,
    inout wire D2DS_X2_Y3,
    inout wire D2DS_X2_Y4,
    inout wire D2DS_X2_Y5,
    inout wire D2DS_X3_Y2,
    inout wire D2DS_X3_Y3,
    inout wire D2DS_X3_Y4,
    inout wire D2DS_X3_Y5,
    inout wire D2DS_X9_Y1,
    inout wire D2DS_X10_Y1,
    inout wire D2DS_X2_Y1,
    inout wire D2DS_X4_Y1,
    inout wire D2DS_X4_Y2,
    inout wire D2DS_X4_Y3,
    inout wire D2DS_X3_Y1,
    inout wire D2DS_X5_Y1,
    inout wire D2DS_X5_Y4,
    inout wire D2DS_X5_Y5,
    inout wire D2DS_X7_Y1,
    inout wire D2DS_X6_Y2,
    inout wire D2DS_X5_Y2,
    inout wire D2DS_X6_Y4,
    inout wire D2DS_X8_Y1,
    inout wire D2DS_X6_Y1,
    inout wire D2DS_X6_Y3,
    inout wire D2DS_X6_Y5,
    inout wire D2DS_X4_Y4,
    inout wire D2DS_X4_Y5,
    inout wire D2DS_X5_Y3,
    inout wire D2DW_X0_Y10,
    inout wire D2DW_X0_Y9,
    inout wire D2DW_X0_Y8,
    inout wire D2DW_X0_Y7,
    inout wire D2DW_X0_Y6,
    inout wire D2DW_X0_Y5,
    inout wire D2DW_X0_Y4,
    inout wire D2DW_X0_Y3,
    inout wire D2DW_X0_Y2,
    inout wire D2DW_X0_Y1,
    inout wire D2DW_X0_Y0,
    inout wire D2DW_X5_Y8,
    inout wire D2DW_X5_Y7,
    inout wire D2DW_X5_Y6,
    inout wire D2DW_X4_Y6,
    inout wire D2DW_X3_Y6,
    inout wire D2DW_X2_Y6,
    inout wire D2DW_X1_Y6,
    inout wire D2DW_X5_Y5,
    inout wire D2DW_X4_Y5,
    inout wire D2DW_X3_Y5,
    inout wire D2DW_X2_Y5,
    inout wire D2DW_X5_Y4,
    inout wire D2DW_X4_Y4,
    inout wire D2DW_X3_Y4,
    inout wire D2DW_X2_Y4,
    inout wire D2DW_X5_Y3,
    inout wire D2DW_X5_Y2,
    inout wire D2DW_X5_Y1,
    inout wire D2DW_X1_Y4,
    inout wire D2DW_X1_Y5,
    inout wire D2DW_X5_Y0,
    inout wire D2DW_X1_Y0,
    inout wire D2DW_X1_Y1,
    inout wire D2DW_X1_Y2,
    inout wire D2DW_X1_Y3,
    inout wire D2DW_X2_Y0,
    inout wire D2DW_X2_Y1,
    inout wire D2DW_X2_Y2,
    inout wire D2DW_X2_Y3,
    inout wire D2DW_X3_Y0,
    inout wire D2DW_X3_Y1,
    inout wire D2DW_X3_Y2,
    inout wire D2DW_X3_Y3,
    inout wire D2DW_X4_Y0,
    inout wire D2DW_X4_Y1,
    inout wire D2DW_X4_Y2,
    inout wire D2DW_X4_Y3,
    inout wire D2DW_X1_Y7,
    inout wire D2DW_X1_Y8,
    inout wire D2DW_X1_Y9,
    inout wire D2DW_X1_Y10,
    inout wire D2DW_X2_Y7,
    inout wire D2DW_X2_Y8,
    inout wire D2DW_X2_Y9,
    inout wire D2DW_X2_Y10,
    inout wire D2DW_X3_Y7,
    inout wire D2DW_X3_Y8,
    inout wire D2DW_X3_Y9,
    inout wire D2DW_X3_Y10,
    inout wire D2DW_X4_Y7,
    inout wire D2DW_X4_Y8,
    inout wire D2DW_X4_Y9,
    inout wire D2DW_X4_Y10,
    inout wire D2DW_X5_Y10,
    inout wire D2DW_X5_Y9
);

  hemaia i_hemaia (
      .io_clk_i(CRTL_X1_Y3),
      .io_rst_ni(CRTL_X1_Y1),
      .io_bypass_pll_division_i(CRTL_X1_Y4),
      .io_clk_obs_o(CRBL_X5_Y2),
      .io_clk_periph_i(CRTL_X2_Y4),
      .io_rst_periph_ni(CRTL_X1_Y0),
      .io_test_mode_i(CRTL_X1_Y2),
      .io_chip_id_i({
        CRBL_X2_Y1,
        CRBL_X3_Y1,
        CRBL_X4_Y1,
        CRBL_X5_Y1,
        CRBR_X0_Y1,
        CRBR_X1_Y1,
        CRBR_X2_Y1,
        CRBR_X3_Y1
      }),
      .io_boot_mode_i(CRBL_X3_Y4),
      .io_east_test_being_requested_i(CRTR_X3_Y0),
      .io_east_test_request_o(CRTR_X2_Y1),
      .io_flow_control_east_rts_o(CRBR_X2_Y4),
      .io_flow_control_east_cts_i(CRBR_X2_Y5),
      .io_flow_control_east_rts_i(CRBR_X2_Y3),
      .io_flow_control_east_cts_o(CRBR_X1_Y3),
      .io_east_d2d({
        D2DE_X3_Y10,
        D2DE_X3_Y9,
        D2DE_X3_Y8,
        D2DE_X3_Y7,
        D2DE_X2_Y10,
        D2DE_X2_Y9,
        D2DE_X2_Y8,
        D2DE_X2_Y7,
        D2DE_X1_Y10,
        D2DE_X1_Y9,
        D2DE_X1_Y8,
        D2DE_X1_Y7,
        D2DE_X0_Y10,
        D2DE_X0_Y9,
        D2DE_X0_Y8,
        D2DE_X0_Y7,
        D2DE_X4_Y10,
        D2DE_X4_Y9,
        D2DE_X5_Y9,
        D2DE_X5_Y8,
        D2DE_X4_Y8,
        D2DE_X4_Y7,
        D2DE_X4_Y3,
        D2DE_X4_Y2,
        D2DE_X3_Y6,
        D2DE_X4_Y6,
        D2DE_X4_Y4,
        D2DE_X3_Y4,
        D2DE_X2_Y6,
        D2DE_X4_Y5,
        D2DE_X3_Y5,
        D2DE_X2_Y4,
        D2DE_X1_Y6,
        D2DE_X1_Y5,
        D2DE_X1_Y4,
        D2DE_X0_Y4,
        D2DE_X0_Y6,
        D2DE_X0_Y5,
        D2DE_X5_Y5,
        D2DE_X5_Y4,
        D2DE_X3_Y3,
        D2DE_X3_Y2,
        D2DE_X3_Y1,
        D2DE_X3_Y0,
        D2DE_X2_Y3,
        D2DE_X2_Y2,
        D2DE_X2_Y1,
        D2DE_X2_Y0,
        D2DE_X1_Y3,
        D2DE_X1_Y2,
        D2DE_X1_Y1,
        D2DE_X1_Y0,
        D2DE_X0_Y3,
        D2DE_X0_Y2,
        D2DE_X0_Y1,
        D2DE_X0_Y0,
        D2DE_X4_Y1,
        D2DE_X4_Y0,
        D2DE_X5_Y1,
        D2DE_X5_Y0
      }),
      .io_west_test_being_requested_i(CRTL_X2_Y2),
      .io_west_test_request_o(CRTL_X2_Y3),
      .io_flow_control_west_rts_o(CRBL_X2_Y2),
      .io_flow_control_west_cts_i(CRBL_X2_Y4),
      .io_flow_control_west_rts_i(CRBL_X3_Y3),
      .io_flow_control_west_cts_o(CRBL_X2_Y3),
      .io_west_d2d({
        D2DW_X4_Y10,
        D2DW_X4_Y9,
        D2DW_X4_Y8,
        D2DW_X4_Y7,
        D2DW_X3_Y10,
        D2DW_X3_Y9,
        D2DW_X3_Y8,
        D2DW_X3_Y7,
        D2DW_X2_Y10,
        D2DW_X2_Y9,
        D2DW_X2_Y8,
        D2DW_X2_Y7,
        D2DW_X1_Y10,
        D2DW_X1_Y9,
        D2DW_X1_Y8,
        D2DW_X1_Y7,
        D2DW_X5_Y10,
        D2DW_X5_Y9,
        D2DW_X0_Y10,
        D2DW_X0_Y9,
        D2DW_X5_Y8,
        D2DW_X5_Y7,
        D2DW_X5_Y3,
        D2DW_X5_Y2,
        D2DW_X4_Y6,
        D2DW_X5_Y6,
        D2DW_X5_Y4,
        D2DW_X4_Y4,
        D2DW_X3_Y6,
        D2DW_X5_Y5,
        D2DW_X4_Y5,
        D2DW_X3_Y4,
        D2DW_X2_Y6,
        D2DW_X2_Y5,
        D2DW_X2_Y4,
        D2DW_X1_Y4,
        D2DW_X1_Y6,
        D2DW_X1_Y5,
        D2DW_X0_Y6,
        D2DW_X0_Y5,
        D2DW_X4_Y3,
        D2DW_X4_Y2,
        D2DW_X4_Y1,
        D2DW_X4_Y0,
        D2DW_X3_Y3,
        D2DW_X3_Y2,
        D2DW_X3_Y1,
        D2DW_X3_Y0,
        D2DW_X2_Y3,
        D2DW_X2_Y2,
        D2DW_X2_Y1,
        D2DW_X2_Y0,
        D2DW_X1_Y3,
        D2DW_X1_Y2,
        D2DW_X1_Y1,
        D2DW_X1_Y0,
        D2DW_X5_Y1,
        D2DW_X5_Y0,
        D2DW_X0_Y2,
        D2DW_X0_Y1
      }),
      .io_north_test_being_requested_i(CRTL_X3_Y3),
      .io_north_test_request_o(CRTL_X4_Y3),
      .io_flow_control_north_rts_o(CRTR_X3_Y2),
      .io_flow_control_north_cts_i(CRTR_X0_Y2),
      .io_flow_control_north_rts_i(CRTR_X2_Y2),
      .io_flow_control_north_cts_o(CRTR_X1_Y2),
      .io_north_d2d({
        D2DN_X10_Y4,
        D2DN_X10_Y3,
        D2DN_X10_Y2,
        D2DN_X10_Y1,
        D2DN_X9_Y4,
        D2DN_X9_Y3,
        D2DN_X9_Y2,
        D2DN_X9_Y1,
        D2DN_X8_Y4,
        D2DN_X8_Y3,
        D2DN_X8_Y2,
        D2DN_X8_Y1,
        D2DN_X7_Y4,
        D2DN_X7_Y3,
        D2DN_X7_Y2,
        D2DN_X7_Y1,
        D2DN_X10_Y0,
        D2DN_X9_Y0,
        D2DN_X10_Y5,
        D2DN_X9_Y5,
        D2DN_X6_Y4,
        D2DN_X6_Y2,
        D2DN_X6_Y0,
        D2DN_X8_Y0,
        D2DN_X6_Y3,
        D2DN_X5_Y1,
        D2DN_X6_Y1,
        D2DN_X7_Y0,
        D2DN_X5_Y4,
        D2DN_X5_Y3,
        D2DN_X5_Y0,
        D2DN_X3_Y0,
        D2DN_X4_Y2,
        D2DN_X4_Y1,
        D2DN_X4_Y0,
        D2DN_X2_Y0,
        D2DN_X4_Y4,
        D2DN_X4_Y3,
        D2DN_X6_Y5,
        D2DN_X5_Y5,
        D2DN_X3_Y4,
        D2DN_X3_Y3,
        D2DN_X3_Y2,
        D2DN_X3_Y1,
        D2DN_X2_Y4,
        D2DN_X2_Y3,
        D2DN_X2_Y2,
        D2DN_X2_Y1,
        D2DN_X1_Y4,
        D2DN_X1_Y3,
        D2DN_X1_Y2,
        D2DN_X1_Y1,
        D2DN_X0_Y4,
        D2DN_X0_Y3,
        D2DN_X0_Y2,
        D2DN_X0_Y1,
        D2DN_X1_Y0,
        D2DN_X0_Y0,
        D2DN_X2_Y5,
        D2DN_X1_Y5
      }),
      .io_south_test_being_requested_i(CRBL_X4_Y2),
      .io_south_test_request_o(CRBL_X3_Y2),
      .io_flow_control_south_rts_o(CRBR_X0_Y2),
      .io_flow_control_south_cts_i(CRBR_X2_Y2),
      .io_flow_control_south_rts_i(CRBR_X1_Y2),
      .io_flow_control_south_cts_o(CRBR_X0_Y3),
      .io_south_d2d({
        D2DS_X10_Y5,
        D2DS_X10_Y4,
        D2DS_X10_Y3,
        D2DS_X10_Y2,
        D2DS_X9_Y5,
        D2DS_X9_Y4,
        D2DS_X9_Y3,
        D2DS_X9_Y2,
        D2DS_X8_Y5,
        D2DS_X8_Y4,
        D2DS_X8_Y3,
        D2DS_X8_Y2,
        D2DS_X7_Y5,
        D2DS_X7_Y4,
        D2DS_X7_Y3,
        D2DS_X7_Y2,
        D2DS_X10_Y1,
        D2DS_X9_Y1,
        D2DS_X9_Y0,
        D2DS_X8_Y0,
        D2DS_X6_Y5,
        D2DS_X6_Y3,
        D2DS_X6_Y1,
        D2DS_X8_Y1,
        D2DS_X6_Y4,
        D2DS_X5_Y2,
        D2DS_X6_Y2,
        D2DS_X7_Y1,
        D2DS_X5_Y5,
        D2DS_X5_Y4,
        D2DS_X5_Y1,
        D2DS_X3_Y1,
        D2DS_X4_Y3,
        D2DS_X4_Y2,
        D2DS_X4_Y1,
        D2DS_X2_Y1,
        D2DS_X4_Y5,
        D2DS_X4_Y4,
        D2DS_X5_Y0,
        D2DS_X4_Y0,
        D2DS_X3_Y5,
        D2DS_X3_Y4,
        D2DS_X3_Y3,
        D2DS_X3_Y2,
        D2DS_X2_Y5,
        D2DS_X2_Y4,
        D2DS_X2_Y3,
        D2DS_X2_Y2,
        D2DS_X1_Y5,
        D2DS_X1_Y4,
        D2DS_X1_Y3,
        D2DS_X1_Y2,
        D2DS_X0_Y5,
        D2DS_X0_Y4,
        D2DS_X0_Y3,
        D2DS_X0_Y2,
        D2DS_X1_Y1,
        D2DS_X0_Y1,
        D2DS_X1_Y0,
        D2DS_X0_Y0
      }),
      .io_uart_tx_o(CRBL_X1_Y4),
      .io_uart_rx_i(CRBL_X1_Y3),
      .io_uart_rts_no(CRBL_X1_Y2),
      .io_uart_cts_ni(CRBL_X1_Y1),
      .io_gpio({CRBR_X3_Y2, CRBR_X3_Y3, CRBR_X3_Y4, CRBR_X3_Y5}),
      .io_spim_sck_o(CRTL_X3_Y4),
      .io_spim_csb_o(CRTL_X4_Y4),
      .io_spim_sd({CRTR_X3_Y3, CRTR_X2_Y3, CRTR_X1_Y3, CRTR_X0_Y3}),
      .io_i2c_sda(CRTL_X2_Y1),
      .io_i2c_scl(CRTL_X2_Y0),
      .io_jtag_trst_ni(CRTR_X4_Y3),
      .io_jtag_tck_i(CRTR_X4_Y2),
      .io_jtag_tms_i(CRTR_X4_Y1),
      .io_jtag_tdi_i(CRTR_X4_Y0),
      .io_jtag_tdo_o(CRTR_X3_Y1)
  );
endmodule
