
/* This alias module is for use internal to the netlister only.
 Please
     do not use the same name for modules or
 assume the existence of 
    this module. */

module cds_alias (
    cds_alias_sig,
    cds_alias_sig
);

  parameter width = 1;

  input [width:1] cds_alias_sig;

endmodule
